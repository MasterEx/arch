-- Ntanasis Periklis A.M.:3070130 - Xatzipetros Mixail A.M.:3070175
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY regfile IS
GENERIC (
n : INTEGER := 16
);
PORT (
Write1				: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
Clock, Write1AD 	: IN STD_LOGIC;
Read1AD, Read2AD	: IN STD_LOGIC;
Read1, Read2		: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0)
Output				: OUT STD_LOGIC_VECTOR((8*n)-1 DOWNTO 0)
);
END regfile;


ARCHITECTURE behavior OF regfile IS

--SIGNAL Output :	STD_LOGIC_VECTOR(n-1 DOWNTO 0);
COMPONENT reg
PORT (
D 		: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
Resetn 	: IN STD_LOGIC;
E, Clock: IN STD_LOGIC;
Q 		: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0)
);
END COMPONENT;

COMPONENT reg0
PORT (
D 		: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
Resetn 	: IN STD_LOGIC;
E, Clock: IN STD_LOGIC;
Q 		: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0)
);
END COMPONENT;

BEGIN
	PROCESS (Clock)
	BEGIN
		
	END PROCESS;
END behavior;
